//-------------------------------------------------------------------------
//      VGA controller                                                   --
//      Kyle Kloepper                                                    --
//      4-05-2005                                                        --
//                                                                       --
//      Modified by Stephen Kempf 04-08-2005                             --
//                                10-05-2006                             --
//                                03-12-2007                             --
//      Translated by Joe Meng    07-07-2013                             --
//      Modified by Po-Han Huang  12-08-2017                             --
//      Spring 2018 Distribution                                         --
//                                                                       --
//      Used standard 640x480 vga found at epanorama                     --
//                                                                       --
//      reference: http://www.xilinx.com/bvdocs/userguides/ug130.pdf     --
//                 http://www.epanorama.net/documents/pc/vga_timing.html --
//                                                                       --
//      note: The standard is changed slightly because of 25 mhz instead --
//            of 25.175 mhz pixel clock. Refresh rate drops slightly.    --
//                                                                       --
//      For use with ECE 385 Lab 8 and Final Project                     --
//      ECE Department @ UIUC                                            --
//-------------------------------------------------------------------------

/**
 * Module: vga_controller
 * Input: clk, reset, vga_clk
 * Output: vga_hs, vga_vs, vga_blank_n, vga_sync_n, [9:0] vga_x, [9:0] vga_y
 * Description: This module handle VGA timming and generate VGA control 
                signals. It also outputs current VGA pixel coordinates for
                other control routines.
 */

module  vga_controller (input              clk,         // 50 MHz clock
                                           reset,       // Active-high reset signal
                        output logic       vga_hs,      // Horizontal sync pulse.  Active low
                                           vga_vs,      // Vertical sync pulse.  Active low
                        input              vga_clk,     // 25 MHz VGA clock input
                        output logic       vga_blank_n, // Blanking interval indicator.  Active low.
                                           vga_sync_n,  // Composite Sync signal.  Active low.  We don't use it in this lab,
                                                        //     but the video DAC on the DE2 board requires an input for it.
                        output logic [9:0] vga_x,      // horizontal coordinate
                                           vga_y       // vertical coordinate
                        );     
    
    // 800 pixels per line (including front/back porch)
    // 525 lines per frame (including front/back porch)
    parameter [9:0] H_TOTAL = 10'd800;
    parameter [9:0] V_TOTAL = 10'd525;
    
    logic vga_hs_in, vga_vs_in, vga_blank_n_in;
    logic [9:0] h_counter, v_counter;
    logic [9:0] h_counter_in, v_counter_in;
    
    assign vga_sync_n = 1'b0;
    assign vga_x = h_counter;
    assign vga_y = v_counter;
    
    // VGA control signals. 
    // vga_clk is generated by PLL, so you will have to manually generate it in simulation.
    always_ff @ (posedge vga_clk)
    begin
        if (reset)
        begin
            vga_hs <= 1'b0;
            vga_vs <= 1'b0;
            vga_blank_n <= 1'b0;
            h_counter <= 10'd0;
            v_counter <= 10'd0;
        end
        else
        begin
            vga_hs <= vga_hs_in;
            vga_vs <= vga_vs_in;
            vga_blank_n <= vga_blank_n_in;
            h_counter <= h_counter_in;
            v_counter <= v_counter_in;
        end
    end
    
    always_comb
    begin
        // Horizontal and vertical counter
        h_counter_in = h_counter + 10'd1;
        v_counter_in = v_counter;
        if (h_counter + 10'd1 == H_TOTAL)
        begin
            h_counter_in = 10'd0;
            if (v_counter + 10'd1 == V_TOTAL) v_counter_in = 10'd0;
            else v_counter_in = v_counter + 10'd1;
        end
        // Horizontal sync pulse is 96 pixels long at pixels 656-752
        // (Signal is registered to ensure clean output waveform)
        vga_hs_in = 1'b1;
        if (h_counter_in >= 10'd656 && h_counter_in < 10'd752) vga_hs_in = 1'b0;

        // Vertical sync pulse is 2 lines (800 pixels each) long at line 490-491
        // (Signal is registered to ensure clean output waveform)
        vga_vs_in = 1'b1;
        if (v_counter_in >= 10'd490 && v_counter_in < 10'd492) vga_vs_in = 1'b0;

        // Display pixels (inhibit blanking) between horizontal 0-639 and vertical 0-479 (640x480)
        vga_blank_n_in = 1'b0;
        if (h_counter_in < 10'd640 && v_counter_in < 10'd480) vga_blank_n_in = 1'b1;
    end
    
endmodule
